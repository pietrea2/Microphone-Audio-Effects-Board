��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��$�����Q�-E�zW�l5n$�0��4WO�G&z��|��T�<��r��Xz�q�*���*i�В-L_O�B��pL����V����d��Gc]%��u���c��D����gP�������������44��Pg��w�k�n�L�t�=�ʠ̲J�=�	�$tG�讧��p,��sC��Xu�_ S�	��mZK�qnu�*u"ǋ<�L*�2S���!��i�އh���
������)�=k��l��hx��I��} ���l��CaoK^G����F�HE���}�-���8���C��)�6v��q+���BɃ״��0�Ўl���Ax�`93Di�j�]��0x��uHo8ȁ�h�+���]�,L��uS��|�>5��9�8>�U̒ �|�o=���{�
'�[	��ԄgI.��Rs���Z�GݲB�_/h�_g�ˢGmYAa/E���,Ӥ`�΁b�d�@��+
��kz<ˤ(�w����0C݊��L87�C��������z��H�w��ڻJ�:>A��>I�B	�KW�-H��
 �ѶJ��;�\�16Ji�,�z}�:d�9E��_����Z���o-�[Ɯ��F$v�KG�%Z�:�oA4w�)[����:��z�X�o=B�e|�_2��ͰUSo����I#ظu��#x	oC}�v�%����KBU�2 p3 e�+�0ʝ��l�;$랉�A��t�h�?\�<��d"]���xuB�@3�{��e40/���GC��������ھΛ�HWR4��M�q��q��x�Gf�5�AW@{�-��LX�d��փ��Z�$�|�t��u�z(t�]7C�ua�Q�t��>l̘�9qaD���5:Ee��LsQ���荌'�^��[`xXP���-�����欜y��������nl�U��s#��{�&�@�%*�A#l2��HQr�Z�w���h�a+@Wfp��Md��S��#��uQMĹ)�8���^�J%+3�i�����1�J-��S+��h�ۼ�%�d�FP[ �Z�+]#�*
B���ĭӔt]���Vg��J)�_?Ir^lD�����3e�ݬ�.���J�?����j,=u�PH��<T^�.�,x��Ҭ�}�M�x���#��ed䋩�+�?R-W��g-4Hsć@-�O����$U��k�)�2��f�6�Ūۚ��3���=����,�-L��(��MS�D�b~v�9H��w^c�\���a$|�������ө�}4�^ԥ �0���$�/�@�Q
�Y2}Rp��rRu�8\�JݢCUсp�l�Y��4�IVKĺN����5K��S����U�<��$!%����4
��\�O��&��?�pI����|�b>�7�m>\8H�������Y��ǒa,��J�����������)�aR�rqp�ޤ.K����e�pҜ�>M���m�	|����x�q��C5̗�ދ\oa��<][ݨW������m}'3&_���+	V0��K���o7]��L���k�S�~�� ��Kݕՙ�N�$�&�ǂ��M�
���u���zR#=�%�n mEIq�w���!:���6[�U-���P}��k*EAd�x�D�帷,�N����N�����xb�P[��<%��e��xtRG�D(Q��$6M*����,���=3�k�tcp���\9�%�rO���J/ud�N�!���CRp�z���x�Ӳ�X�S��?T�vTW/�{�OK��~ck��z��ibw�����/�ꮡ�;u�N/����4%s4�a��9\o2�	���ɀ�1�c������\N��)��x�B��Z�2{�\�J@=Z�� Q|�4���6Ӻ蟴8uHߞ�m��\�n���m�F����>�F�����L��￲5ۻ��_��C�+�a�\%G�*�3����s6��D��d�����I�N���d*�1i�|�-�oS��L&�Y~>��%���@���o�-^�8��%<����8�5�}¬&t4ԁOKƊJ�dܫh٫�D��������#Yo��v\�l�����G@C�9�\���ӿ(4`�v�X��zO��C�l&�3
(�%����Ύ7Q�
��9������3��E�(�7����=w�wy��S�Jb��ռ�k��)9
��_J�Q���ޤ�f��|)O����&]<�H'��)���w'x�=P�3�D.'f�I��6�d��"���_ֱA�ș�q�9і}z1>p׽֘,�#G�Z�Ǎ����
0���Rt���Z[%l8bp��kT^љ>9ԆtY<I��f�22���>��o�̄i�v�}����[�`��{u4�5��̂�p��OKdzn'I��"��Ϲ/�0pӨ�1W��>^�q����~��Q�Rj���[i�&�Ua�u @�q\��������B�y��WY�sxK_u|��m�/a�9�Mf��?�����j=��>��
����d��p�Q�e�h�ʭ1���CH��K��0��v����*_AX3���J���A�N�U��b+]YԸA�ݝ������Џ4;�1��c�5������3��_G�Xai�S8��+�y�hq�d��7��nm�����νa:✋��KKl�f�U`��zc��y^�3:�0儘Lp&�Ͼ	)Gd8M�.P�uP�?�#krV��/07(��ÏBN�f�G��������RP��F>��uA^}kl{ڧ���*���~�n�'��B;����F�"mY���p�
Ĥ�]���ܚe؀�lh����K�e�_4�
�(h�|��$-r2��\s�ۤڀ����z�c��qJ�F�b����GA��/���6�����0���4��,��ݳ����$������.K@1+�9��̒��ύ�pG��|��G�Z�[I��)���� F��4ԇ�L�"{{��Һ�dao��n���F/�p�3�(jTW��I��0�I�[�$Q��� s��\�)��봜���C�:M�C\
m6h�q?�<�-�C\����0����H$,q{wT�]Ӵ����>Z���Gݎ���]
��:��yR$���k�`a�|	���%y=u��"~�~{�F"� 4s�G�R����S��{H�Hdx�f8P�Hͤd�g=b`Y��|��`�iQ�n���#��klnӻ�P3�"B�i��#����)����/���HuͲ��Ì���m���N��6�zL	6H�N6;(ed�s(�
u�QUW<�I���P7��C�e$�o{Ü���&:��cё
�!!��!D���<�g^խUn�6�{��B�7���*�J���oR�:��iÃ��5�(�o�,8�x��\��,/Q�}�����h�˩���/�r��Zf� �j@�BIQO .��N��װ�J7� �)|v}㽠�/ȯ����z�
uc�Fyv���i)T��\o��d`\Tq��V� �	uN��~ �6�B� �b~�&�_`���:�o�� ����p��^B�ɜ�dp��G�f�b��Y����58W�����p��������	W�p����r�Om��$<'���a�f��8��������y�r���*#�=V��WACM�A�=��63G�~���^ض��DiBqX ǧ�������H�Y���`_fi��,W^72�M%���>e
[핑�n�B��ESD���Ơ�3��7�A�.Æ�*�!�-��B�2�	�+�0�d��5�iu0u�Sf��\~����H��EL���'�#"�S_����z�Hq_��8[���3�z�������$F�č�6�t��aJ�ӝg_��D���Y������ ��-��AN#��b�SZ �n��Gq�gSV������6+{�=ׯ����@�d���.�Bz����E� ��\+�0���n�.�w��$ת>x�{�һDҴ+�coIN#�q���q�C!���k �< �SlY�:�Dl^@�:{ғ�������2��E���N����~ˏ:��*�w��&!��J�����J�A>�5��U�8�"!���a�Etߵ�i>�4p�B�n`���e'�aʈ�a���X+#�!�+|�}I�)���pm(��ТBCڍn��<I��Q�~Q	���(�E���[8��WL}3��ȩ�g��ߨ����ҧ�����Z�b�߸90MR�?����3���٬�H���₹�@iQ�,���$C��&^���}�x{�a��!�vK)�������Q��΄���C��� �Ĉ�	86l�q���hM��^����#��@y��,
0>���F�l�;]!Q����wk���Z�wư�0���h*��Lno���v��M�q#�T!9&�o��(����E?I�GCF�$�9��B4	] 7�_�t+0r���O�^����Z��Y%���LFN���ckh�7(i��"a�3\e�ǎwl|-NVj�m��n7��NO�5Tg/9�ܣ��r[ZT��)�rTk�S>-��,�;zo;1ʥ0H������?�{ma�����q'�2�)x����GM���y7Z�W����+����k��1�	��e���'���
S��n����*�t~,�M]��&2>Dۛi(*TL��Y��1���t��&�Y�&���3L��o���X��7Y*&H�]��J�kua�@k�,����~I��VȒ��]���U+�I�|RW J0�צ��
�#vW�ݨ����l,���L������+�����p
�S���w��T��,~&6�Lؚ;Nk��#}i~P/#j)�a$h�s�F�rU��)���<�>���mE��Xh�૟�A��_�#�+�Iw:�P�*>^��N�*�o^�N�.�(�������IZ\`V�{�"~������)?��`k$W~�&+� u���z�=���Ȧu�]���8�/�zײ֞����a�o>�⸛��E�k2/����vU{b�w���
��e���H��Z���w��rM����:q����j��뼦[��l��Z��k����Yr�i�l��U���[z�@�s|!����oP���e0ը~��(�!�0�dv�|ߨ9vnn�^��񔼉\
ǭ["ڰ�����zS��DF^�ꕍ]�vޢ��BҚ6�tNbp&*� �R�`��MiU�)������i�a8hfd�c��	:�?�mQ�ٱTk�G������I0`*�Vոl���1��IM߈�	>M9��b�Tl;1���c��	[�6�u����������3 \7(��V/���&��\�ơ�^��2�1n@Ej�V������,����j`��s���)�@��������t'A71���f�H[�W�O8�p,��n�s'N���.bU�8�`.t��fo�m�'ԣ��*�$�ѬEŜ�1��k; ��y	s0�6��1����΅(���#�С�)�"ڤ�7L���d�N_aH���Ƭ��1Χ��c��~Y��僚V>��h�'ɘ���e�@"�$D���G�����3<���o;���6X%5�1/^C{%��qۙe�cl-�q=ģ�I���y�T�N�ۊ���Ԫ���Ͻu���I(�AHb�����yU^M��:,*?n��S����DS��ߊ���̼"��!��~����:>�ȑ2G.�s��|�E�a���a�v(`�d�6&�{�N����%&/��6 �����%'"�����2�i�=S��OR3q�f���䋦��W]'��h~7s6 C�!�*���#>F�>t�0���]���jR�����U dL��%N��v��̯�6�]!�VS��a����܍?Ck�簂nRqw�p4}�YJD-ܩj�����y-���C��ʱ�i�R1{ �=�&F��6QR����xa����[ZFEhHjE%���&H�[��OQ�1��/Ȱ=aϾ���P�m�c7��v�������;[�5��[��]3-�P%_�ծ�U�T�>S�-��!��1�����!���܆�2gsáa*Y�\�T��G��C(��bXR:��4��it�Ұ<W�o;���sƞҧ�*lRě�0GA��?*��C�(2�x���+PN �A��d:KA�F$ ���6A��N���~]�L�hG,#=��63��ʒD�6g�N�`��|R��;o/҉h�����RfB&��!����#�RZ���ZV�j��s^��c2��iʲ�h�.	�]<6Ï�Kw�U��z"K>���=���c�G����^��!n�{�Beڦ*�7w֯w�~������;��\"�=n�fI��4&ڱ���ҷ%ӥ`��,7d�V��G�*X
<���X�4�k����,]�hҒ1d��u$zWt�Q5t��u+�[��i�ںN���Q����v��4A}W�d�y!���v]� ;(}�����ԟ�!���btB�G_Sv�&�#��q�aǝ�`�V)�uc�t_Z;3-���5�_Z�RG�ޅ��S���	���Þ<c���5�,�����4ƙ�ǃ���|��r1�u%5Z&�[�������kV��L��bt�O��P7�En��V#�h\�n):��]�h6�kl�WH&�u1��6�� �76q��P�E��}	y�?e�y���D�,G�4����5|^U��e���J؁ftc�M(_|E�$�}vX�������x2�����ފ/1 ^F��l$
��e�q W'���C	,I�g<=�[�p"��ۼ�ڲ�a����~)5{�?Y_�"W��K�Jn��(Q����z5�v�m  ��~��TT��ԭ��2'�+�R�v�K|��G����wg,�B���#�3�D��͕\���Ȏ\VD��V�?|�[GX"�;��N�`���^S��)
q�Iyr���ٵ�@6��<���9��r���"=�6Z��	�v�B��i�'�ED���ʰx��ı6�Q_����c�$,h���V?���2S# ��,q���i�O��z��m���X�Dͷ���gX��=�#���$��l�h�>חm[�%�aK8�ɕ�awzk<� ��ܿ{4�+=����8��Ρ(G� �a1:�;��խ�mV�[70���^���2��	j'�p�V�S���:~2(��nej+�y�B�(��-fH��eC�HN�X����n�<$�Q�l�;�����p�~��3Ê�9�c
�\�E�'���1���'2��p��
C��M0��65Xjv�0˻��#�|?�XK���_���E<����m�zN5�Gu�W
�v>��Z`�i��Uf8�O�x�X&L��'���!;Ѵ[B�v�J�*�Y�˵G���i���C����0h�E�xΫ���B"@9���ѧ�dZ�ժ����6���Wy��L�y�03�/�Vٚ�̓Bn�"nݾ}VY�-�^eKRtv��B��X�x3��c7#�RnєWDy�4)����Ы�?~�I+��4�
��`��4Z����Xj�t�)���,&��x�g��޺��B�
�%�P�[(�ɏ������'�z����<�q�#�L����o:+�jd��M�%��U%�#'$����v����w�,}�ލ���^��)!P(��)>mLq��S!�jb_��P6)��6�V�Ȳ.bī����ԯ_\�YH<k����;ǤS��S�� ���U
3��� yI��x�'�Z��%G�x���Y�􍻨a���'��CO��E�u��j��V+�gH���*�sw��:�	�����-P�P�� +��f{����C�^�o�� ^����l�����HI�h�r�=G4���C2�Y��S���$٥��a�.�C	���C��t�ߝ)��A� |��幜&Rr�BK~��q����xL���
	���5�|J�o�]a��s�Ԯu�0=�R�*_pHEۜv��-�g@E�T�m��S��y��XT�C�4+�`��}zGd-ᴿ%)��"�B��HG��^h�W�?�N��<���� ��}�
ew��IdK�x`j��*fmI�`��b+�m�W�u�it�� Z2�F	}��?����iךR�2^u���О�-�F�tAM�{�](S΋��>O���®u���܇S��	2��#953�4NɔD�L�j��)�`wi�a3o<�XN�F,���]�uGӾEpt헌��Ի�}@"ڛ4'ӹ�jn9ɸ��FM]�2�-=q�h�/�u�X�;�orBv�K8������$�	+�Hg+�8V_V0A<D��|�p��ؽ��*��2_�0�w~�.��sP1�EYAJ��G��:~Q�CuN�&�j=ML	A� �ٜ��#Ԕ�Ҳ�L�I���Q��6�}}p�ҹ�5�M��	
�>�p��;�v�{�"��-:�h�]<�a��X��N,c������[����sB��x���X�t7w@4S��UW.�3��QEۋ�]�+������9��6�Q����͐5o�'�I�ة�����E��(���=粝qRs��Nl�E8R���~�g)�D��}{N��>�NO�Ĳohz�2B7��j�DI9�k��t�J��Y��	��Z��_|!���Y�^�-�b^V�C�Ǒ΃B���p.�U��5����"��t��ݒ��'�nu95�t��^e� �*����z�>���$�-���9h�����UM;|��zq�\[����W.г������4�SC��۞�?��;��>�k)��\����n���=�~{��� @�$8��ݿeG!a��l�`�����m3:�eo��/�|�!K����1�љ���!�d����8o�2YY�*|�t�;�6�7-�9�w��8TY�lό.*cܝ����:���[k�@>xM�:��Kw�-�jJ���~�%���e���b�W]E�K���QU�}�����d��D6ŝj���΄`� ��q�o�ݓg?�^ ���&�X����ܪ8GG�˾��<豋���N�䄅V%b��4Y�;���k��v/Y 9 ��%����(E��Ax�������$�k��a��?�t@���Tξ�b����f� �s�W�dׇ�5L]/�  �&ѕ��0�|�zW=H�vF��$3� �/`��*D��8�� -��1u��n')dX��z*�����Yd{�z����5L����J3'x0hL���V�.�;:�d>`%���؋��N��<`��H|4l�9^����R�{���=pN�0�m��'�/1���-�9�|��s̉������uË-^N�몮��b�C 8��a��8��e,*[�_j G�3���1���3����7��*�G�s��nd������'��~����fт�_O�����4�+�@���i����P#Vcе*��Y���#Ҵ���xm�!��)'����3U�5U�  ��;�Kp�0�&�㡦�c�ZhߚH�
ػe�HZ6e��mM�O:���L�Fjt.����$Z �?-��#�\EF�WB�`�R\���5Ű���l*��v�Sт��Z1~��O*K�ꖠ�Z�tB��~�y[u�9�)_r(�k��h2��Ƥ��)]��j�0vt�S:��`f��O�ć�1c�$'=m�&�v/����`Q��)Ԝ�>�N%a���HP���1����w���
�ʆO݋ٿݤ��S��x�,g��Ⱦ%�>c3�ۄ>��H��z����/������*kF��8A�Wׅ�R�[��´q��"��j�ǻ"�ڷ�F�ș�ó�[�D�?P&A���GWy���e��	��*L�0�^���/tjq?sH�8�>���}.ka�' �{�)s��L��ܤ!���Z�%�sFT5��?�"0��;��;�&��4����J�@
����M����+�,�l��1����t���ɰWE�	Fv�C��� C?ň�$8���j@PA�j,#wgP��Rh�g[��Ĺ��Ђ�x���b%{_P%~7$W�]k�������)�_(i��s9��=��8���$٪8��>��\+�Y�;���.���}� �'��o��˜h���3Q�E�r��*��Kd~�b�tТf�X��P�2�X�&��+����C��B*(wT�}@��ȝaS���̼���'s�t�Q	�oQ0���(�7�
i�G����H���=��h�ǈH�`LZ�wB���a�?	�_Iu_���;��_�suc��Q�y�����f�|����$[�Bj&�O���Յ�a�y�F��_� ���ط7�����"�2r���fшe��>_W,��1��*��>LY�1���F�H�����2&F�����_l\� ����#s7�tT�qƤK��d�y�r�i�v�op�o�3�,�z9X���RW�`�Asx��)Τ��YN^j� ,Ė�X��1� ާ�!(M�~��؜Z�[�ӧ�%���/)�تcT�5�1�Ќr>�#U�1�5����![H�>���Y&��G���R߰`ۈԐk.����л����Љ��0}�v���c�t�vA����A ��C=nUұ}����4�6������Z�v�.�㙦��������٨�L�@��0�4��.fF�:c@L�zyg��o�:�0�[�J����u�BXka$ȦY�r��#�Q�DZ��!�L���C��|�ڮ���S��0x·ت�	e�)J�2��d �Z����~�+ZX9T7^�د�HD���D�?"r{S̛B��Z���i�/�@��o=_'�ڑ���ͺ�7݄X�P��z�/-�
���>?ǌ[)
����η���@����������·w\��T�d�sUf�;�a���Q�O�����r^C��[���%��nj��Rj�}��oy��Vw����>rm۪��T@j�Oʵ��\~��!�Q]��p{��a��|�.���4�f�s��Z���G[��Z�a�����Y/	�3��L��J�gS����S��f 1���o#m��[�|߻�i�Vp���N�y��FS��WԛJ&�p+�̶���&�_M���I%�ݱ-J�w���b���̣-��u	ͽ���^C+9������X,󮸀��Fȡ���(�lD��z�����)����[*9 [�t� s�)�F����ږ�?��E����|%J\R.�<[FYVJ��JxmS�jWdK`cB����Ǔ�'q�<��#�Nވ�#=1s"HҥR���K�6-����7�z�ÿ�}�#^U:´>�[���ضndE�`#�>d�p����s/�h�R�VnՋeU�c���G���X�u�����ken��4��u��xIJm��574�1�w���r@Mča� �����9�܌��%��cρב�hvJ���������Ue����ú3�Ru&��yl*��w�4,��A:�YV�l��C�K��A0�-�T�ƙ�X˽���K�"����3 f+��b��#�ݿ��E�/޲��X� ���䇳&�~,PMs��	̋"4Sr��_~I;:SVڷ������8r��B�M�ӽ�|��OPz�2���4�s����y�f;�r�!�ؖ�D.���?Avi�I��?��ڣ��"����t�fz����&eeӳli�{�p ���t1�U�˶	uo������Ž�$��s:�W���8��d+�\޿�1<�{��Jxx]����c.�P�?W��*1[����c��$uc�I0�^���_>��U�kI�{�i����\v��m:f�^���6����֪���Hd�E��A]Wq�������)W�.E:�д����>L�������[9���9d-��5���HꊽZ�Z���m�R�٭�kM-<�_Dl=kM)���~s�]����:�Ʒe�
�ut7�ɺ8�|�tP-x����mLB�Jx6.WD������论L-;%�5d�8v�MɃ�缿�����i��Z/��@�t������,k�㧬�I�Z���z>�������I�5�[p�L��(��1��7O ��O�{y*@{�ҥ��}�̐d�I���m?q��T�2�a���Ȇ�Ea�L��E�2��XD�,�l:ݹ �dp����]��ý�Γ�Hd��:i�]�4��n��K��'���-��*��xQ��^g��-�d�l'�X�VZ�|��,[%�ĥ�Kc!,Q Io���.&�k�WҦ���r^�����$���G�ytM��9���1x�� &�	{�WLq��yU{c�W!��